library IEEE;
use ieee.std_logic_1164.all;
use ieee.STD_LOGIC_UNSIGNED.all;
use std.textio.all;
use work.aux_functions.all;

entity RAM_mem is
      
end RAM_mem;

architecture RAM_mem of RAM_mem is 
begin

end RAM_mem;