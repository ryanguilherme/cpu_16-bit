library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity register_file_tb is
	-- Port ();
end register_file_tb;

architecture Behavorial 
